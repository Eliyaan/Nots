module main

@[inline]
fn ceil(nb f64) int {
	return -int(-nb)
}