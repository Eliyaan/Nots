
module main

struct Junction {
mut:
	destroyed bool
	in_gate   bool
	x         i64
	y         i64
}